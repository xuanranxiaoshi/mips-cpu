`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/01/04 20:55:51
// Design Name: 
// Module Name: tb_inst_mem_dual
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 测试双端口指令ROM的可行性
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_inst_mem_dual();
    reg clk;
    reg rst;
    
endmodule
