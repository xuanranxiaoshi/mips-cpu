// decode 是否访存
`define MEM_LOAD 2'b01
`define MEM_STOR 2'b10
`define MEM_NOT 2'b00 //not mem instruction